
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
--use work.ALU_components_pack.all;

entity bin_to_bcd_lut8 is
   port ( 
			binary_in : in  unsigned(7 downto 0);  -- binary input width
			bcd_out   : out std_logic_vector(9 downto 0)   -- BCD output, 10 bits [2|4|4] to display a 3 digit BCD value when input has length 8
		);
end bin_to_bcd_lut8;

architecture structural of bin_to_bcd_lut8 is 

begin  
	-- DEVELOPE YOUR CODE HERE
	process (binary_in)
	begin
		case binary_in is
           when "00000000" => bcd_out <= "0000000000";
            when "00000001" => bcd_out <= "0000000001";
            when "00000010" => bcd_out <= "0000000010";
            when "00000011" => bcd_out <= "0000000011";
            when "00000100" => bcd_out <= "0000000100";
            when "00000101" => bcd_out <= "0000000101";
            when "00000110" => bcd_out <= "0000000110";
            when "00000111" => bcd_out <= "0000000111";
            when "00001000" => bcd_out <= "0000001000";
            when "00001001" => bcd_out <= "0000001001";
            when "00001010" => bcd_out <= "0000010000";
            when "00001011" => bcd_out <= "0000010001";
            when "00001100" => bcd_out <= "0000010010";
            when "00001101" => bcd_out <= "0000010011";
            when "00001110" => bcd_out <= "0000010100";
            when "00001111" => bcd_out <= "0000010101";
            when "00010000" => bcd_out <= "0000010110";
            when "00010001" => bcd_out <= "0000010111";
            when "00010010" => bcd_out <= "0000011000";
            when "00010011" => bcd_out <= "0000011001";
            when "00010100" => bcd_out <= "0000100000";
            when "00010101" => bcd_out <= "0000100001";
            when "00010110" => bcd_out <= "0000100010";
            when "00010111" => bcd_out <= "0000100011";
            when "00011000" => bcd_out <= "0000100100";
            when "00011001" => bcd_out <= "0000100101";
            when "00011010" => bcd_out <= "0000100110";
            when "00011011" => bcd_out <= "0000100111";
            when "00011100" => bcd_out <= "0000101000";
            when "00011101" => bcd_out <= "0000101001";
            when "00011110" => bcd_out <= "0000110000";
            when "00011111" => bcd_out <= "0000110001";
            when "00100000" => bcd_out <= "0000110010";
            when "00100001" => bcd_out <= "0000110011";
            when "00100010" => bcd_out <= "0000110100";
            when "00100011" => bcd_out <= "0000110101";
            when "00100100" => bcd_out <= "0000110110";
            when "00100101" => bcd_out <= "0000110111";
            when "00100110" => bcd_out <= "0000111000";
            when "00100111" => bcd_out <= "0000111001";
            when "00101000" => bcd_out <= "0001000000";
            when "00101001" => bcd_out <= "0001000001";
            when "00101010" => bcd_out <= "0001000010";
            when "00101011" => bcd_out <= "0001000011";
            when "00101100" => bcd_out <= "0001000100";
            when "00101101" => bcd_out <= "0001000101";
            when "00101110" => bcd_out <= "0001000110";
            when "00101111" => bcd_out <= "0001000111";
            when "00110000" => bcd_out <= "0001001000";
            when "00110001" => bcd_out <= "0001001001";
            when "00110010" => bcd_out <= "0001010000";
            when "00110011" => bcd_out <= "0001010001";
            when "00110100" => bcd_out <= "0001010010";
            when "00110101" => bcd_out <= "0001010011";
            when "00110110" => bcd_out <= "0001010100";
            when "00110111" => bcd_out <= "0001010101";
            when "00111000" => bcd_out <= "0001010110";
            when "00111001" => bcd_out <= "0001010111";
            when "00111010" => bcd_out <= "0001011000";
            when "00111011" => bcd_out <= "0001011001";
            when "00111100" => bcd_out <= "0001100000";
            when "00111101" => bcd_out <= "0001100001";
            when "00111110" => bcd_out <= "0001100010";
            when "00111111" => bcd_out <= "0001100011";
            when "01000000" => bcd_out <= "0001100100";
            when "01000001" => bcd_out <= "0001100101";
            when "01000010" => bcd_out <= "0001100110";
            when "01000011" => bcd_out <= "0001100111";
            when "01000100" => bcd_out <= "0001101000";
            when "01000101" => bcd_out <= "0001101001";
            when "01000110" => bcd_out <= "0001110000";
            when "01000111" => bcd_out <= "0001110001";
            when "01001000" => bcd_out <= "0001110010";
            when "01001001" => bcd_out <= "0001110011";
            when "01001010" => bcd_out <= "0001110100";
            when "01001011" => bcd_out <= "0001110101";
            when "01001100" => bcd_out <= "0001110110";
            when "01001101" => bcd_out <= "0001110111";
            when "01001110" => bcd_out <= "0001111000";
            when "01001111" => bcd_out <= "0001111001";
            when "01010000" => bcd_out <= "0010000000";
            when "01010001" => bcd_out <= "0010000001";
            when "01010010" => bcd_out <= "0010000010";
            when "01010011" => bcd_out <= "0010000011";
            when "01010100" => bcd_out <= "0010000100";
            when "01010101" => bcd_out <= "0010000101";
            when "01010110" => bcd_out <= "0010000110";
            when "01010111" => bcd_out <= "0010000111";
            when "01011000" => bcd_out <= "0010001000";
            when "01011001" => bcd_out <= "0010001001";
            when "01011010" => bcd_out <= "0010010000";
            when "01011011" => bcd_out <= "0010010001";
            when "01011100" => bcd_out <= "0010010010";
            when "01011101" => bcd_out <= "0010010011";
            when "01011110" => bcd_out <= "0010010100";
            when "01011111" => bcd_out <= "0010010101";
            when "01100000" => bcd_out <= "0010010110";
            when "01100001" => bcd_out <= "0010010111";
            when "01100010" => bcd_out <= "0010011000";
            when "01100011" => bcd_out <= "0010011001";
            when "01100100" => bcd_out <= "0100000000";
            when "01100101" => bcd_out <= "0100000001";
            when "01100110" => bcd_out <= "0100000010";
            when "01100111" => bcd_out <= "0100000011";
            when "01101000" => bcd_out <= "0100000100";
            when "01101001" => bcd_out <= "0100000101";
            when "01101010" => bcd_out <= "0100000110";
            when "01101011" => bcd_out <= "0100000111";
            when "01101100" => bcd_out <= "0100001000";
            when "01101101" => bcd_out <= "0100001001";
            when "01101110" => bcd_out <= "0100010000";
            when "01101111" => bcd_out <= "0100010001";
            when "01110000" => bcd_out <= "0100010010";
            when "01110001" => bcd_out <= "0100010011";
            when "01110010" => bcd_out <= "0100010100";
            when "01110011" => bcd_out <= "0100010101";
            when "01110100" => bcd_out <= "0100010110";
            when "01110101" => bcd_out <= "0100010111";
            when "01110110" => bcd_out <= "0100011000";
            when "01110111" => bcd_out <= "0100011001";
            when "01111000" => bcd_out <= "0100100000";
            when "01111001" => bcd_out <= "0100100001";
            when "01111010" => bcd_out <= "0100100010";
            when "01111011" => bcd_out <= "0100100011";
            when "01111100" => bcd_out <= "0100100100";
            when "01111101" => bcd_out <= "0100100101";
            when "01111110" => bcd_out <= "0100100110";
            when "01111111" => bcd_out <= "0100100111";
            when "10000000" => bcd_out <= "0100101000";
            when "10000001" => bcd_out <= "0100101001";
            when "10000010" => bcd_out <= "0100110000";
            when "10000011" => bcd_out <= "0100110001";
            when "10000100" => bcd_out <= "0100110010";
            when "10000101" => bcd_out <= "0100110011";
            when "10000110" => bcd_out <= "0100110100";
            when "10000111" => bcd_out <= "0100110101";
            when "10001000" => bcd_out <= "0100110110";
            when "10001001" => bcd_out <= "0100110111";
            when "10001010" => bcd_out <= "0100111000";
            when "10001011" => bcd_out <= "0100111001";
            when "10001100" => bcd_out <= "0101000000";
            when "10001101" => bcd_out <= "0101000001";
            when "10001110" => bcd_out <= "0101000010";
            when "10001111" => bcd_out <= "0101000011";
            when "10010000" => bcd_out <= "0101000100";
            when "10010001" => bcd_out <= "0101000101";
            when "10010010" => bcd_out <= "0101000110";
            when "10010011" => bcd_out <= "0101000111";
            when "10010100" => bcd_out <= "0101001000";
            when "10010101" => bcd_out <= "0101001001";
            when "10010110" => bcd_out <= "0101010000";
            when "10010111" => bcd_out <= "0101010001";
            when "10011000" => bcd_out <= "0101010010";
            when "10011001" => bcd_out <= "0101010011";
            when "10011010" => bcd_out <= "0101010100";
            when "10011011" => bcd_out <= "0101010101";
            when "10011100" => bcd_out <= "0101010110";
            when "10011101" => bcd_out <= "0101010111";
            when "10011110" => bcd_out <= "0101011000";
            when "10011111" => bcd_out <= "0101011001";
            when "10100000" => bcd_out <= "0101100000";
            when "10100001" => bcd_out <= "0101100001";
            when "10100010" => bcd_out <= "0101100010";
            when "10100011" => bcd_out <= "0101100011";
            when "10100100" => bcd_out <= "0101100100";
            when "10100101" => bcd_out <= "0101100101";
            when "10100110" => bcd_out <= "0101100110";
            when "10100111" => bcd_out <= "0101100111";
            when "10101000" => bcd_out <= "0101101000";
            when "10101001" => bcd_out <= "0101101001";
            when "10101010" => bcd_out <= "0101110000";
            when "10101011" => bcd_out <= "0101110001";
            when "10101100" => bcd_out <= "0101110010";
            when "10101101" => bcd_out <= "0101110011";
            when "10101110" => bcd_out <= "0101110100";
            when "10101111" => bcd_out <= "0101110101";
            when "10110000" => bcd_out <= "0101110110";
            when "10110001" => bcd_out <= "0101110111";
            when "10110010" => bcd_out <= "0101111000";
            when "10110011" => bcd_out <= "0101111001";
            when "10110100" => bcd_out <= "0110000000";
            when "10110101" => bcd_out <= "0110000001";
            when "10110110" => bcd_out <= "0110000010";
            when "10110111" => bcd_out <= "0110000011";
            when "10111000" => bcd_out <= "0110000100";
            when "10111001" => bcd_out <= "0110000101";
            when "10111010" => bcd_out <= "0110000110";
            when "10111011" => bcd_out <= "0110000111";
            when "10111100" => bcd_out <= "0110001000";
            when "10111101" => bcd_out <= "0110001001";
            when "10111110" => bcd_out <= "0110010000";
            when "10111111" => bcd_out <= "0110010001";
            when "11000000" => bcd_out <= "0110010010";
            when "11000001" => bcd_out <= "0110010011";
            when "11000010" => bcd_out <= "0110010100";
            when "11000011" => bcd_out <= "0110010101";
            when "11000100" => bcd_out <= "0110010110";
            when "11000101" => bcd_out <= "0110010111";
            when "11000110" => bcd_out <= "0110011000";
            when "11000111" => bcd_out <= "0110011001";
            when "11001000" => bcd_out <= "1000000000";
            when "11001001" => bcd_out <= "1000000001";
            when "11001010" => bcd_out <= "1000000010";
            when "11001011" => bcd_out <= "1000000011";
            when "11001100" => bcd_out <= "1000000100";
            when "11001101" => bcd_out <= "1000000101";
            when "11001110" => bcd_out <= "1000000110";
            when "11001111" => bcd_out <= "1000000111";
            when "11010000" => bcd_out <= "1000001000";
            when "11010001" => bcd_out <= "1000001001";
            when "11010010" => bcd_out <= "1000010000";
            when "11010011" => bcd_out <= "1000010001";
            when "11010100" => bcd_out <= "1000010010";
            when "11010101" => bcd_out <= "1000010011";
            when "11010110" => bcd_out <= "1000010100";
            when "11010111" => bcd_out <= "1000010101";
            when "11011000" => bcd_out <= "1000010110";
            when "11011001" => bcd_out <= "1000010111";
            when "11011010" => bcd_out <= "1000011000";
            when "11011011" => bcd_out <= "1000011001";
            when "11011100" => bcd_out <= "1000100000";
            when "11011101" => bcd_out <= "1000100001";
            when "11011110" => bcd_out <= "1000100010";
            when "11011111" => bcd_out <= "1000100011";
            when "11100000" => bcd_out <= "1000100100";
            when "11100001" => bcd_out <= "1000100101";
            when "11100010" => bcd_out <= "1000100110";
            when "11100011" => bcd_out <= "1000100111";
            when "11100100" => bcd_out <= "1000101000";
            when "11100101" => bcd_out <= "1000101001";
            when "11100110" => bcd_out <= "1000110000";
            when "11100111" => bcd_out <= "1000110001";
            when "11101000" => bcd_out <= "1000110010";
            when "11101001" => bcd_out <= "1000110011";
            when "11101010" => bcd_out <= "1000110100";
            when "11101011" => bcd_out <= "1000110101";
            when "11101100" => bcd_out <= "1000110110";
            when "11101101" => bcd_out <= "1000110111";
            when "11101110" => bcd_out <= "1000111000";
            when "11101111" => bcd_out <= "1000111001";
            when "11110000" => bcd_out <= "1001000000";
            when "11110001" => bcd_out <= "1001000001";
            when "11110010" => bcd_out <= "1001000010";
            when "11110011" => bcd_out <= "1001000011";
            when "11110100" => bcd_out <= "1001000100";
            when "11110101" => bcd_out <= "1001000101";
            when "11110110" => bcd_out <= "1001000110";
            when "11110111" => bcd_out <= "1001000111";
            when "11111000" => bcd_out <= "1001001000";
            when "11111001" => bcd_out <= "1001001001";
            when "11111010" => bcd_out <= "1001010000";
            when "11111011" => bcd_out <= "1001010001";
            when "11111100" => bcd_out <= "1001010010";
            when "11111101" => bcd_out <= "1001010011";
            when "11111110" => bcd_out <= "1001010100";
            when "11111111" => bcd_out <= "1001010101";
 
			when others => null;
		end case;
	end process;
end structural;
		
	