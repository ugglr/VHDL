
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
--use work.ALU_components_pack.all;

entity bin_to_bcd_lut10 is
   port ( 
			binary_in : in  unsigned(9 downto 0);  -- binary input width
			bcd_out   : out std_logic_vector(11 downto 0)   -- BCD output, 10 bits [2|4|4] to display a 3 digit BCD value when input has length 8
		);
end bin_to_bcd_lut10;

architecture structural of bin_to_bcd_lut10 is 

begin  
	-- DEVELOPE YOUR CODE HERE
	process (binary_in)
	begin
		case binary_in is           when "0000000000" => bcd_out <= "000000000000"; --0
            when "0000000001" => bcd_out <= "000000000001"; --001
            when "0000000010" => bcd_out <= "000000000010"; --002
            when "0000000011" => bcd_out <= "000000000011"; --003
            when "0000000100" => bcd_out <= "000000000100"; --004
            when "0000000101" => bcd_out <= "000000000101"; --005
            when "0000000110" => bcd_out <= "000000000110"; --006
            when "0000000111" => bcd_out <= "000000000111"; --007
            when "0000001000" => bcd_out <= "000000001000"; --008
            when "0000001001" => bcd_out <= "000000001001"; --009
            when "0000001010" => bcd_out <= "000000000001"; --01
            when "0000001011" => bcd_out <= "000000010001"; --011
            when "0000001100" => bcd_out <= "000000010010"; --012
            when "0000001101" => bcd_out <= "000000010011"; --013
            when "0000001110" => bcd_out <= "000000010100"; --014
            when "0000001111" => bcd_out <= "000000010101"; --015
            when "0000010000" => bcd_out <= "000000010110"; --016
            when "0000010001" => bcd_out <= "000000010111"; --017
            when "0000010010" => bcd_out <= "000000011000"; --018
            when "0000010011" => bcd_out <= "000000011001"; --019
            when "0000010100" => bcd_out <= "000000000010"; --02
            when "0000010101" => bcd_out <= "000000100001"; --021
            when "0000010110" => bcd_out <= "000000100001"; --021
            when "0000010111" => bcd_out <= "000000100010"; --022
            when "0000011000" => bcd_out <= "000000100011"; --023
            when "0000011001" => bcd_out <= "000000100100"; --024
            when "0000011010" => bcd_out <= "000000100101"; --025
            when "0000011011" => bcd_out <= "000000100110"; --026
            when "0000011100" => bcd_out <= "000000100111"; --027
            when "0000011101" => bcd_out <= "000000101000"; --028
            when "0000011110" => bcd_out <= "000000101001"; --029
            when "0000011111" => bcd_out <= "000000000011"; --03
            when "0000100000" => bcd_out <= "000000110001"; --031
            when "0000100001" => bcd_out <= "000000110010"; --032
            when "0000100010" => bcd_out <= "000000110011"; --033
            when "0000100011" => bcd_out <= "000000110100"; --034
            when "0000100100" => bcd_out <= "000000110101"; --035
            when "0000100101" => bcd_out <= "000000110110"; --036
            when "0000100110" => bcd_out <= "000000110111"; --037
            when "0000100111" => bcd_out <= "000000111000"; --038
            when "0000101000" => bcd_out <= "000000111001"; --039
            when "0000101001" => bcd_out <= "000000000100"; --04
            when "0000101010" => bcd_out <= "000001000001"; --041
            when "0000101011" => bcd_out <= "000001000010"; --042
            when "0000101100" => bcd_out <= "000001000011"; --043
            when "0000101101" => bcd_out <= "000001000100"; --044
            when "0000101110" => bcd_out <= "000001000101"; --045
            when "0000101111" => bcd_out <= "000001000110"; --046
            when "0000110000" => bcd_out <= "000001000111"; --047
            when "0000110001" => bcd_out <= "000001001000"; --048
            when "0000110010" => bcd_out <= "000001001001"; --049
            when "0000110011" => bcd_out <= "000000000101"; --05
            when "0000110100" => bcd_out <= "000001010001"; --051
            when "0000110101" => bcd_out <= "000001010010"; --052
            when "0000110110" => bcd_out <= "000001010011"; --053
            when "0000110111" => bcd_out <= "000001010100"; --054
            when "0000111000" => bcd_out <= "000001010101"; --055
            when "0000111001" => bcd_out <= "000001010110"; --056
            when "0000111010" => bcd_out <= "000001010111"; --057
            when "0000111011" => bcd_out <= "000001011000"; --058
            when "0000111100" => bcd_out <= "000001011001"; --059
            when "0000111101" => bcd_out <= "000000000110"; --06
            when "0000111110" => bcd_out <= "000001100001"; --061
            when "0000111111" => bcd_out <= "000001100010"; --062
            when "0001000000" => bcd_out <= "000001100011"; --063
            when "0001000001" => bcd_out <= "000001100011"; --063
            when "0001000010" => bcd_out <= "000001100100"; --064
            when "0001000011" => bcd_out <= "000001100101"; --065
            when "0001000100" => bcd_out <= "000001100110"; --066
            when "0001000101" => bcd_out <= "000001100111"; --067
            when "0001000110" => bcd_out <= "000001101000"; --068
            when "0001000111" => bcd_out <= "000001101001"; --069
            when "0001001000" => bcd_out <= "000000000111"; --07
            when "0001001001" => bcd_out <= "000001110001"; --071
            when "0001001010" => bcd_out <= "000001110010"; --072
            when "0001001011" => bcd_out <= "000001110011"; --073
            when "0001001100" => bcd_out <= "000001110100"; --074
            when "0001001101" => bcd_out <= "000001110101"; --075
            when "0001001110" => bcd_out <= "000001110110"; --076
            when "0001001111" => bcd_out <= "000001110111"; --077
            when "0001010000" => bcd_out <= "000001111000"; --078
            when "0001010001" => bcd_out <= "000001111001"; --079
            when "0001010010" => bcd_out <= "000000001000"; --08
            when "0001010011" => bcd_out <= "000010000001"; --081
            when "0001010100" => bcd_out <= "000010000010"; --082
            when "0001010101" => bcd_out <= "000010000011"; --083
            when "0001010110" => bcd_out <= "000010000100"; --084
            when "0001010111" => bcd_out <= "000010000101"; --085
            when "0001011000" => bcd_out <= "000010000110"; --086
            when "0001011001" => bcd_out <= "000010000111"; --087
            when "0001011010" => bcd_out <= "000010001000"; --088
            when "0001011011" => bcd_out <= "000010001001"; --089
            when "0001011100" => bcd_out <= "000000001001"; --09
            when "0001011101" => bcd_out <= "000010010001"; --091
            when "0001011110" => bcd_out <= "000010010010"; --092
            when "0001011111" => bcd_out <= "000010010011"; --093
            when "0001100000" => bcd_out <= "000010010100"; --094
            when "0001100001" => bcd_out <= "000010010101"; --095
            when "0001100010" => bcd_out <= "000010010110"; --096
            when "0001100011" => bcd_out <= "000010010111"; --097
            when "0001100100" => bcd_out <= "000010011000"; --098
            when "0001100101" => bcd_out <= "000010011001"; --099
            when "0001100110" => bcd_out <= "000000000001"; --1
            when "0001100111" => bcd_out <= "000100000001"; --101
            when "0001101000" => bcd_out <= "000100000010"; --102
            when "0001101001" => bcd_out <= "000100000011"; --103
            when "0001101010" => bcd_out <= "000100000100"; --104
            when "0001101011" => bcd_out <= "000100000100"; --104
            when "0001101100" => bcd_out <= "000100000101"; --105
            when "0001101101" => bcd_out <= "000100000110"; --106
            when "0001101110" => bcd_out <= "000100000111"; --107
            when "0001101111" => bcd_out <= "000100001000"; --108
            when "0001110000" => bcd_out <= "000100001001"; --109
            when "0001110001" => bcd_out <= "000000010001"; --11
            when "0001110010" => bcd_out <= "000100010001"; --111
            when "0001110011" => bcd_out <= "000100010010"; --112
            when "0001110100" => bcd_out <= "000100010011"; --113
            when "0001110101" => bcd_out <= "000100010100"; --114
            when "0001110110" => bcd_out <= "000100010101"; --115
            when "0001110111" => bcd_out <= "000100010110"; --116
            when "0001111000" => bcd_out <= "000100010111"; --117
            when "0001111001" => bcd_out <= "000100011000"; --118
            when "0001111010" => bcd_out <= "000100011001"; --119
            when "0001111011" => bcd_out <= "000000010010"; --12
            when "0001111100" => bcd_out <= "000100100001"; --121
            when "0001111101" => bcd_out <= "000100100010"; --122
            when "0001111110" => bcd_out <= "000100100011"; --123
            when "0001111111" => bcd_out <= "000100100100"; --124
            when "0010000000" => bcd_out <= "000100100101"; --125
            when "0010000001" => bcd_out <= "000100100110"; --126
            when "0010000010" => bcd_out <= "000100100111"; --127
            when "0010000011" => bcd_out <= "000100101000"; --128
            when "0010000100" => bcd_out <= "000100101001"; --129
            when "0010000101" => bcd_out <= "000000010011"; --13
            when "0010000110" => bcd_out <= "000100110001"; --131
            when "0010000111" => bcd_out <= "000100110010"; --132
            when "0010001000" => bcd_out <= "000100110011"; --133
            when "0010001001" => bcd_out <= "000100110100"; --134
            when "0010001010" => bcd_out <= "000100110101"; --135
            when "0010001011" => bcd_out <= "000100110110"; --136
            when "0010001100" => bcd_out <= "000100110111"; --137
            when "0010001101" => bcd_out <= "000100111000"; --138
            when "0010001110" => bcd_out <= "000100111001"; --139
            when "0010001111" => bcd_out <= "000000010100"; --14
            when "0010010000" => bcd_out <= "000101000001"; --141
            when "0010010001" => bcd_out <= "000101000010"; --142
            when "0010010010" => bcd_out <= "000101000011"; --143
            when "0010010011" => bcd_out <= "000101000100"; --144
            when "0010010100" => bcd_out <= "000101000101"; --145
            when "0010010101" => bcd_out <= "000101000110"; --146
            when "0010010110" => bcd_out <= "000101000110"; --146
            when "0010010111" => bcd_out <= "000101000111"; --147
            when "0010011000" => bcd_out <= "000101001000"; --148
            when "0010011001" => bcd_out <= "000101001001"; --149
            when "0010011010" => bcd_out <= "000000010101"; --15
            when "0010011011" => bcd_out <= "000101010001"; --151
            when "0010011100" => bcd_out <= "000101010010"; --152
            when "0010011101" => bcd_out <= "000101010011"; --153
            when "0010011110" => bcd_out <= "000101010100"; --154
            when "0010011111" => bcd_out <= "000101010101"; --155
            when "0010100000" => bcd_out <= "000101010110"; --156
            when "0010100001" => bcd_out <= "000101010111"; --157
            when "0010100010" => bcd_out <= "000101011000"; --158
            when "0010100011" => bcd_out <= "000101011001"; --159
            when "0010100100" => bcd_out <= "000000010110"; --16
            when "0010100101" => bcd_out <= "000101100001"; --161
            when "0010100110" => bcd_out <= "000101100010"; --162
            when "0010100111" => bcd_out <= "000101100011"; --163
            when "0010101000" => bcd_out <= "000101100100"; --164
            when "0010101001" => bcd_out <= "000101100101"; --165
            when "0010101010" => bcd_out <= "000101100110"; --166
            when "0010101011" => bcd_out <= "000101100111"; --167
            when "0010101100" => bcd_out <= "000101101000"; --168
            when "0010101101" => bcd_out <= "000101101001"; --169
            when "0010101110" => bcd_out <= "000000010111"; --17
            when "0010101111" => bcd_out <= "000101110001"; --171
            when "0010110000" => bcd_out <= "000101110010"; --172
            when "0010110001" => bcd_out <= "000101110011"; --173
            when "0010110010" => bcd_out <= "000101110100"; --174
            when "0010110011" => bcd_out <= "000101110101"; --175
            when "0010110100" => bcd_out <= "000101110110"; --176
            when "0010110101" => bcd_out <= "000101110111"; --177
            when "0010110110" => bcd_out <= "000101111000"; --178
            when "0010110111" => bcd_out <= "000101111001"; --179
            when "0010111000" => bcd_out <= "000000011000"; --18
            when "0010111001" => bcd_out <= "000110000001"; --181
            when "0010111010" => bcd_out <= "000110000010"; --182
            when "0010111011" => bcd_out <= "000110000011"; --183
            when "0010111100" => bcd_out <= "000110000100"; --184
            when "0010111101" => bcd_out <= "000110000101"; --185
            when "0010111110" => bcd_out <= "000110000110"; --186
            when "0010111111" => bcd_out <= "000110000111"; --187
            when "0011000000" => bcd_out <= "000110001000"; --188
            when "0011000001" => bcd_out <= "000110001000"; --188
            when "0011000010" => bcd_out <= "000110001001"; --189
            when "0011000011" => bcd_out <= "000000011001"; --19
            when "0011000100" => bcd_out <= "000110010001"; --191
            when "0011000101" => bcd_out <= "000110010010"; --192
            when "0011000110" => bcd_out <= "000110010011"; --193
            when "0011000111" => bcd_out <= "000110010100"; --194
            when "0011001000" => bcd_out <= "000110010101"; --195
            when "0011001001" => bcd_out <= "000110010110"; --196
            when "0011001010" => bcd_out <= "000110010111"; --197
            when "0011001011" => bcd_out <= "000110011000"; --198
            when "0011001100" => bcd_out <= "000110011001"; --199
            when "0011001101" => bcd_out <= "000000000010"; --2
            when "0011001110" => bcd_out <= "001000000001"; --201
            when "0011001111" => bcd_out <= "001000000010"; --202
            when "0011010000" => bcd_out <= "001000000011"; --203
            when "0011010001" => bcd_out <= "001000000100"; --204
            when "0011010010" => bcd_out <= "001000000101"; --205
            when "0011010011" => bcd_out <= "001000000110"; --206
            when "0011010100" => bcd_out <= "001000000111"; --207
            when "0011010101" => bcd_out <= "001000001000"; --208
            when "0011010110" => bcd_out <= "001000001001"; --209
            when "0011010111" => bcd_out <= "000000100001"; --21
            when "0011011000" => bcd_out <= "001000010001"; --211
            when "0011011001" => bcd_out <= "001000010010"; --212
            when "0011011010" => bcd_out <= "001000010011"; --213
            when "0011011011" => bcd_out <= "001000010100"; --214
            when "0011011100" => bcd_out <= "001000010101"; --215
            when "0011011101" => bcd_out <= "001000010110"; --216
            when "0011011110" => bcd_out <= "001000010111"; --217
            when "0011011111" => bcd_out <= "001000011000"; --218
            when "0011100000" => bcd_out <= "001000011001"; --219
            when "0011100001" => bcd_out <= "000000100010"; --22
            when "0011100010" => bcd_out <= "001000100001"; --221
            when "0011100011" => bcd_out <= "001000100010"; --222
            when "0011100100" => bcd_out <= "001000100011"; --223
            when "0011100101" => bcd_out <= "001000100100"; --224
            when "0011100110" => bcd_out <= "001000100101"; --225
            when "0011100111" => bcd_out <= "001000100110"; --226
            when "0011101000" => bcd_out <= "001000100111"; --227
            when "0011101001" => bcd_out <= "001000101000"; --228
            when "0011101010" => bcd_out <= "001000101001"; --229
            when "0011101011" => bcd_out <= "001000101001"; --229
            when "0011101100" => bcd_out <= "000000100011"; --23
            when "0011101101" => bcd_out <= "001000110001"; --231
            when "0011101110" => bcd_out <= "001000110010"; --232
            when "0011101111" => bcd_out <= "001000110011"; --233
            when "0011110000" => bcd_out <= "001000110100"; --234
            when "0011110001" => bcd_out <= "001000110101"; --235
            when "0011110010" => bcd_out <= "001000110110"; --236
            when "0011110011" => bcd_out <= "001000110111"; --237
            when "0011110100" => bcd_out <= "001000111000"; --238
            when "0011110101" => bcd_out <= "001000111001"; --239
            when "0011110110" => bcd_out <= "000000100100"; --24
            when "0011110111" => bcd_out <= "001001000001"; --241
            when "0011111000" => bcd_out <= "001001000010"; --242
            when "0011111001" => bcd_out <= "001001000011"; --243
            when "0011111010" => bcd_out <= "001001000100"; --244
            when "0011111011" => bcd_out <= "001001000101"; --245
            when "0011111100" => bcd_out <= "001001000110"; --246
            when "0011111101" => bcd_out <= "001001000111"; --247
            when "0011111110" => bcd_out <= "001001001000"; --248
            when "0011111111" => bcd_out <= "001001001001"; --249
            when "0100000000" => bcd_out <= "000000100101"; --25
            when "0100000001" => bcd_out <= "001001010001"; --251
            when "0100000010" => bcd_out <= "001001010010"; --252
            when "0100000011" => bcd_out <= "001001010011"; --253
            when "0100000100" => bcd_out <= "001001010100"; --254
            when "0100000101" => bcd_out <= "001001010101"; --255
            when "0100000110" => bcd_out <= "001001010110"; --256
            when "0100000111" => bcd_out <= "001001010111"; --257
            when "0100001000" => bcd_out <= "001001011000"; --258
            when "0100001001" => bcd_out <= "001001011001"; --259
            when "0100001010" => bcd_out <= "000000100110"; --26
            when "0100001011" => bcd_out <= "001001100001"; --261
            when "0100001100" => bcd_out <= "001001100010"; --262
            when "0100001101" => bcd_out <= "001001100011"; --263
            when "0100001110" => bcd_out <= "001001100100"; --264
            when "0100001111" => bcd_out <= "001001100101"; --265
            when "0100010000" => bcd_out <= "001001100110"; --266
            when "0100010001" => bcd_out <= "001001100111"; --267
            when "0100010010" => bcd_out <= "001001101000"; --268
            when "0100010011" => bcd_out <= "001001101001"; --269
            when "0100010100" => bcd_out <= "000000100111"; --27
            when "0100010101" => bcd_out <= "001001110001"; --271
            when "0100010110" => bcd_out <= "001001110001"; --271
            when "0100010111" => bcd_out <= "001001110010"; --272
            when "0100011000" => bcd_out <= "001001110011"; --273
            when "0100011001" => bcd_out <= "001001110100"; --274
            when "0100011010" => bcd_out <= "001001110101"; --275
            when "0100011011" => bcd_out <= "001001110110"; --276
            when "0100011100" => bcd_out <= "001001110111"; --277
            when "0100011101" => bcd_out <= "001001111000"; --278
            when "0100011110" => bcd_out <= "001001111001"; --279
            when "0100011111" => bcd_out <= "000000101000"; --28
            when "0100100000" => bcd_out <= "001010000001"; --281
            when "0100100001" => bcd_out <= "001010000010"; --282
            when "0100100010" => bcd_out <= "001010000011"; --283
            when "0100100011" => bcd_out <= "001010000100"; --284
            when "0100100100" => bcd_out <= "001010000101"; --285
            when "0100100101" => bcd_out <= "001010000110"; --286
            when "0100100110" => bcd_out <= "001010000111"; --287
            when "0100100111" => bcd_out <= "001010001000"; --288
            when "0100101000" => bcd_out <= "001010001001"; --289
            when "0100101001" => bcd_out <= "000000101001"; --29
            when "0100101010" => bcd_out <= "001010010001"; --291
            when "0100101011" => bcd_out <= "001010010010"; --292
            when "0100101100" => bcd_out <= "001010010011"; --293
            when "0100101101" => bcd_out <= "001010010100"; --294
            when "0100101110" => bcd_out <= "001010010101"; --295
            when "0100101111" => bcd_out <= "001010010110"; --296
            when "0100110000" => bcd_out <= "001010010111"; --297
            when "0100110001" => bcd_out <= "001010011000"; --298
            when "0100110010" => bcd_out <= "001010011001"; --299
            when "0100110011" => bcd_out <= "000000000011"; --3
            when "0100110100" => bcd_out <= "001100000001"; --301
            when "0100110101" => bcd_out <= "001100000010"; --302
            when "0100110110" => bcd_out <= "001100000011"; --303
            when "0100110111" => bcd_out <= "001100000100"; --304
            when "0100111000" => bcd_out <= "001100000101"; --305
            when "0100111001" => bcd_out <= "001100000110"; --306
            when "0100111010" => bcd_out <= "001100000111"; --307
            when "0100111011" => bcd_out <= "001100001000"; --308
            when "0100111100" => bcd_out <= "001100001001"; --309
            when "0100111101" => bcd_out <= "000000110001"; --31
            when "0100111110" => bcd_out <= "001100010001"; --311
            when "0100111111" => bcd_out <= "001100010010"; --312
            when "0101000000" => bcd_out <= "001100010011"; --313
            when "0101000001" => bcd_out <= "001100010011"; --313
            when "0101000010" => bcd_out <= "001100010100"; --314
            when "0101000011" => bcd_out <= "001100010101"; --315
            when "0101000100" => bcd_out <= "001100010110"; --316
            when "0101000101" => bcd_out <= "001100010111"; --317
            when "0101000110" => bcd_out <= "001100011000"; --318
            when "0101000111" => bcd_out <= "001100011001"; --319
            when "0101001000" => bcd_out <= "000000110010"; --32
            when "0101001001" => bcd_out <= "001100100001"; --321
            when "0101001010" => bcd_out <= "001100100010"; --322
            when "0101001011" => bcd_out <= "001100100011"; --323
            when "0101001100" => bcd_out <= "001100100100"; --324
            when "0101001101" => bcd_out <= "001100100101"; --325
            when "0101001110" => bcd_out <= "001100100110"; --326
            when "0101001111" => bcd_out <= "001100100111"; --327
            when "0101010000" => bcd_out <= "001100101000"; --328
            when "0101010001" => bcd_out <= "001100101001"; --329
            when "0101010010" => bcd_out <= "000000110011"; --33
            when "0101010011" => bcd_out <= "001100110001"; --331
            when "0101010100" => bcd_out <= "001100110010"; --332
            when "0101010101" => bcd_out <= "001100110011"; --333
            when "0101010110" => bcd_out <= "001100110100"; --334
            when "0101010111" => bcd_out <= "001100110101"; --335
            when "0101011000" => bcd_out <= "001100110110"; --336
            when "0101011001" => bcd_out <= "001100110111"; --337
            when "0101011010" => bcd_out <= "001100111000"; --338
            when "0101011011" => bcd_out <= "001100111001"; --339
            when "0101011100" => bcd_out <= "000000110100"; --34
            when "0101011101" => bcd_out <= "001101000001"; --341
            when "0101011110" => bcd_out <= "001101000010"; --342
            when "0101011111" => bcd_out <= "001101000011"; --343
            when "0101100000" => bcd_out <= "001101000100"; --344
            when "0101100001" => bcd_out <= "001101000101"; --345
            when "0101100010" => bcd_out <= "001101000110"; --346
            when "0101100011" => bcd_out <= "001101000111"; --347
            when "0101100100" => bcd_out <= "001101001000"; --348
            when "0101100101" => bcd_out <= "001101001001"; --349
            when "0101100110" => bcd_out <= "000000110101"; --35
            when "0101100111" => bcd_out <= "001101010001"; --351
            when "0101101000" => bcd_out <= "001101010010"; --352
            when "0101101001" => bcd_out <= "001101010011"; --353
            when "0101101010" => bcd_out <= "001101010100"; --354
            when "0101101011" => bcd_out <= "001101010100"; --354
            when "0101101100" => bcd_out <= "001101010101"; --355
            when "0101101101" => bcd_out <= "001101010110"; --356
            when "0101101110" => bcd_out <= "001101010111"; --357
            when "0101101111" => bcd_out <= "001101011000"; --358
            when "0101110000" => bcd_out <= "001101011001"; --359
            when "0101110001" => bcd_out <= "000000110110"; --36
            when "0101110010" => bcd_out <= "001101100001"; --361
            when "0101110011" => bcd_out <= "001101100010"; --362
            when "0101110100" => bcd_out <= "001101100011"; --363
            when "0101110101" => bcd_out <= "001101100100"; --364
            when "0101110110" => bcd_out <= "001101100101"; --365
            when "0101110111" => bcd_out <= "001101100110"; --366
            when "0101111000" => bcd_out <= "001101100111"; --367
            when "0101111001" => bcd_out <= "001101101000"; --368
            when "0101111010" => bcd_out <= "001101101001"; --369
            when "0101111011" => bcd_out <= "000000110111"; --37
            when "0101111100" => bcd_out <= "001101110001"; --371
            when "0101111101" => bcd_out <= "001101110010"; --372
            when "0101111110" => bcd_out <= "001101110011"; --373
            when "0101111111" => bcd_out <= "001101110100"; --374
            when "0110000000" => bcd_out <= "001101110101"; --375
            when "0110000001" => bcd_out <= "001101110110"; --376
            when "0110000010" => bcd_out <= "001101110111"; --377
            when "0110000011" => bcd_out <= "001101111000"; --378
            when "0110000100" => bcd_out <= "001101111001"; --379
            when "0110000101" => bcd_out <= "000000111000"; --38
            when "0110000110" => bcd_out <= "001110000001"; --381
            when "0110000111" => bcd_out <= "001110000010"; --382
            when "0110001000" => bcd_out <= "001110000011"; --383
            when "0110001001" => bcd_out <= "001110000100"; --384
            when "0110001010" => bcd_out <= "001110000101"; --385
            when "0110001011" => bcd_out <= "001110000110"; --386
            when "0110001100" => bcd_out <= "001110000111"; --387
            when "0110001101" => bcd_out <= "001110001000"; --388
            when "0110001110" => bcd_out <= "001110001001"; --389
            when "0110001111" => bcd_out <= "000000111001"; --39
            when "0110010000" => bcd_out <= "001110010001"; --391
            when "0110010001" => bcd_out <= "001110010010"; --392
            when "0110010010" => bcd_out <= "001110010011"; --393
            when "0110010011" => bcd_out <= "001110010100"; --394
            when "0110010100" => bcd_out <= "001110010101"; --395
            when "0110010101" => bcd_out <= "001110010110"; --396
            when "0110010110" => bcd_out <= "001110010110"; --396
            when "0110010111" => bcd_out <= "001110010111"; --397
            when "0110011000" => bcd_out <= "001110011000"; --398
            when "0110011001" => bcd_out <= "001110011001"; --399
            when "0110011010" => bcd_out <= "000000000100"; --4
            when "0110011011" => bcd_out <= "010000000001"; --401
            when "0110011100" => bcd_out <= "010000000010"; --402
            when "0110011101" => bcd_out <= "010000000011"; --403
            when "0110011110" => bcd_out <= "010000000100"; --404
            when "0110011111" => bcd_out <= "010000000101"; --405
            when "0110100000" => bcd_out <= "010000000110"; --406
            when "0110100001" => bcd_out <= "010000000111"; --407
            when "0110100010" => bcd_out <= "010000001000"; --408
            when "0110100011" => bcd_out <= "010000001001"; --409
            when "0110100100" => bcd_out <= "000001000001"; --41
            when "0110100101" => bcd_out <= "010000010001"; --411
            when "0110100110" => bcd_out <= "010000010010"; --412
            when "0110100111" => bcd_out <= "010000010011"; --413
            when "0110101000" => bcd_out <= "010000010100"; --414
            when "0110101001" => bcd_out <= "010000010101"; --415
            when "0110101010" => bcd_out <= "010000010110"; --416
            when "0110101011" => bcd_out <= "010000010111"; --417
            when "0110101100" => bcd_out <= "010000011000"; --418
            when "0110101101" => bcd_out <= "010000011001"; --419
            when "0110101110" => bcd_out <= "000001000010"; --42
            when "0110101111" => bcd_out <= "010000100001"; --421
            when "0110110000" => bcd_out <= "010000100010"; --422
            when "0110110001" => bcd_out <= "010000100011"; --423
            when "0110110010" => bcd_out <= "010000100100"; --424
            when "0110110011" => bcd_out <= "010000100101"; --425
            when "0110110100" => bcd_out <= "010000100110"; --426
            when "0110110101" => bcd_out <= "010000100111"; --427
            when "0110110110" => bcd_out <= "010000101000"; --428
            when "0110110111" => bcd_out <= "010000101001"; --429
            when "0110111000" => bcd_out <= "000001000011"; --43
            when "0110111001" => bcd_out <= "010000110001"; --431
            when "0110111010" => bcd_out <= "010000110010"; --432
            when "0110111011" => bcd_out <= "010000110011"; --433
            when "0110111100" => bcd_out <= "010000110100"; --434
            when "0110111101" => bcd_out <= "010000110101"; --435
            when "0110111110" => bcd_out <= "010000110110"; --436
            when "0110111111" => bcd_out <= "010000110111"; --437
            when "0111000000" => bcd_out <= "010000111000"; --438
            when "0111000001" => bcd_out <= "010000111000"; --438
            when "0111000010" => bcd_out <= "010000111001"; --439
            when "0111000011" => bcd_out <= "000001000100"; --44
            when "0111000100" => bcd_out <= "010001000001"; --441
            when "0111000101" => bcd_out <= "010001000010"; --442
            when "0111000110" => bcd_out <= "010001000011"; --443
            when "0111000111" => bcd_out <= "010001000100"; --444
            when "0111001000" => bcd_out <= "010001000101"; --445
            when "0111001001" => bcd_out <= "010001000110"; --446
            when "0111001010" => bcd_out <= "010001000111"; --447
            when "0111001011" => bcd_out <= "010001001000"; --448
            when "0111001100" => bcd_out <= "010001001001"; --449
            when "0111001101" => bcd_out <= "000001000101"; --45
            when "0111001110" => bcd_out <= "010001010001"; --451
            when "0111001111" => bcd_out <= "010001010010"; --452
            when "0111010000" => bcd_out <= "010001010011"; --453
            when "0111010001" => bcd_out <= "010001010100"; --454
            when "0111010010" => bcd_out <= "010001010101"; --455
            when "0111010011" => bcd_out <= "010001010110"; --456
            when "0111010100" => bcd_out <= "010001010111"; --457
            when "0111010101" => bcd_out <= "010001011000"; --458
            when "0111010110" => bcd_out <= "010001011001"; --459
            when "0111010111" => bcd_out <= "000001000110"; --46
            when "0111011000" => bcd_out <= "010001100001"; --461
            when "0111011001" => bcd_out <= "010001100010"; --462
            when "0111011010" => bcd_out <= "010001100011"; --463
            when "0111011011" => bcd_out <= "010001100100"; --464
            when "0111011100" => bcd_out <= "010001100101"; --465
            when "0111011101" => bcd_out <= "010001100110"; --466
            when "0111011110" => bcd_out <= "010001100111"; --467
            when "0111011111" => bcd_out <= "010001101000"; --468
            when "0111100000" => bcd_out <= "010001101001"; --469
            when "0111100001" => bcd_out <= "000001000111"; --47
            when "0111100010" => bcd_out <= "010001110001"; --471
            when "0111100011" => bcd_out <= "010001110010"; --472
            when "0111100100" => bcd_out <= "010001110011"; --473
            when "0111100101" => bcd_out <= "010001110100"; --474
            when "0111100110" => bcd_out <= "010001110101"; --475
            when "0111100111" => bcd_out <= "010001110110"; --476
            when "0111101000" => bcd_out <= "010001110111"; --477
            when "0111101001" => bcd_out <= "010001111000"; --478
            when "0111101010" => bcd_out <= "010001111001"; --479
            when "0111101011" => bcd_out <= "010001111001"; --479
            when "0111101100" => bcd_out <= "000001001000"; --48
            when "0111101101" => bcd_out <= "010010000001"; --481
            when "0111101110" => bcd_out <= "010010000010"; --482
            when "0111101111" => bcd_out <= "010010000011"; --483
            when "0111110000" => bcd_out <= "010010000100"; --484
            when "0111110001" => bcd_out <= "010010000101"; --485
            when "0111110010" => bcd_out <= "010010000110"; --486
            when "0111110011" => bcd_out <= "010010000111"; --487
            when "0111110100" => bcd_out <= "010010001000"; --488
            when "0111110101" => bcd_out <= "010010001001"; --489
            when "0111110110" => bcd_out <= "000001001001"; --49
            when "0111110111" => bcd_out <= "010010010001"; --491
            when "0111111000" => bcd_out <= "010010010010"; --492
            when "0111111001" => bcd_out <= "010010010011"; --493
            when "0111111010" => bcd_out <= "010010010100"; --494
            when "0111111011" => bcd_out <= "010010010101"; --495
            when "0111111100" => bcd_out <= "010010010110"; --496
            when "0111111101" => bcd_out <= "010010010111"; --497
            when "0111111110" => bcd_out <= "010010011000"; --498
            when "0111111111" => bcd_out <= "010010011001"; --499
            when "1000000000" => bcd_out <= "000000000101"; --5
            when "1000000001" => bcd_out <= "010100000001"; --501
            when "1000000010" => bcd_out <= "010100000010"; --502
            when "1000000011" => bcd_out <= "010100000011"; --503
            when "1000000100" => bcd_out <= "010100000100"; --504
            when "1000000101" => bcd_out <= "010100000101"; --505
            when "1000000110" => bcd_out <= "010100000110"; --506
            when "1000000111" => bcd_out <= "010100000111"; --507
            when "1000001000" => bcd_out <= "010100001000"; --508
            when "1000001001" => bcd_out <= "010100001001"; --509
            when "1000001010" => bcd_out <= "000001010001"; --51
            when "1000001011" => bcd_out <= "010100010001"; --511
            when "1000001100" => bcd_out <= "010100010010"; --512
            when "1000001101" => bcd_out <= "010100010011"; --513
            when "1000001110" => bcd_out <= "010100010100"; --514
            when "1000001111" => bcd_out <= "010100010101"; --515
            when "1000010000" => bcd_out <= "010100010110"; --516
            when "1000010001" => bcd_out <= "010100010111"; --517
            when "1000010010" => bcd_out <= "010100011000"; --518
            when "1000010011" => bcd_out <= "010100011001"; --519
            when "1000010100" => bcd_out <= "000001010010"; --52
            when "1000010101" => bcd_out <= "010100100001"; --521
            when "1000010110" => bcd_out <= "010100100001"; --521
            when "1000010111" => bcd_out <= "010100100010"; --522
            when "1000011000" => bcd_out <= "010100100011"; --523
            when "1000011001" => bcd_out <= "010100100100"; --524
            when "1000011010" => bcd_out <= "010100100101"; --525
            when "1000011011" => bcd_out <= "010100100110"; --526
            when "1000011100" => bcd_out <= "010100100111"; --527
            when "1000011101" => bcd_out <= "010100101000"; --528
            when "1000011110" => bcd_out <= "010100101001"; --529
            when "1000011111" => bcd_out <= "000001010011"; --53
            when "1000100000" => bcd_out <= "010100110001"; --531
            when "1000100001" => bcd_out <= "010100110010"; --532
            when "1000100010" => bcd_out <= "010100110011"; --533
            when "1000100011" => bcd_out <= "010100110100"; --534
            when "1000100100" => bcd_out <= "010100110101"; --535
            when "1000100101" => bcd_out <= "010100110110"; --536
            when "1000100110" => bcd_out <= "010100110111"; --537
            when "1000100111" => bcd_out <= "010100111000"; --538
            when "1000101000" => bcd_out <= "010100111001"; --539
            when "1000101001" => bcd_out <= "000001010100"; --54
            when "1000101010" => bcd_out <= "010101000001"; --541
            when "1000101011" => bcd_out <= "010101000010"; --542
            when "1000101100" => bcd_out <= "010101000011"; --543
            when "1000101101" => bcd_out <= "010101000100"; --544
            when "1000101110" => bcd_out <= "010101000101"; --545
            when "1000101111" => bcd_out <= "010101000110"; --546
            when "1000110000" => bcd_out <= "010101000111"; --547
            when "1000110001" => bcd_out <= "010101001000"; --548
            when "1000110010" => bcd_out <= "010101001001"; --549
            when "1000110011" => bcd_out <= "000001010101"; --55
            when "1000110100" => bcd_out <= "010101010001"; --551
            when "1000110101" => bcd_out <= "010101010010"; --552
            when "1000110110" => bcd_out <= "010101010011"; --553
            when "1000110111" => bcd_out <= "010101010100"; --554
            when "1000111000" => bcd_out <= "010101010101"; --555
            when "1000111001" => bcd_out <= "010101010110"; --556
            when "1000111010" => bcd_out <= "010101010111"; --557
            when "1000111011" => bcd_out <= "010101011000"; --558
            when "1000111100" => bcd_out <= "010101011001"; --559
            when "1000111101" => bcd_out <= "000001010110"; --56
            when "1000111110" => bcd_out <= "010101100001"; --561
            when "1000111111" => bcd_out <= "010101100010"; --562
            when "1001000000" => bcd_out <= "010101100011"; --563
            when "1001000001" => bcd_out <= "010101100011"; --563
            when "1001000010" => bcd_out <= "010101100100"; --564
            when "1001000011" => bcd_out <= "010101100101"; --565
            when "1001000100" => bcd_out <= "010101100110"; --566
            when "1001000101" => bcd_out <= "010101100111"; --567
            when "1001000110" => bcd_out <= "010101101000"; --568
            when "1001000111" => bcd_out <= "010101101001"; --569
            when "1001001000" => bcd_out <= "000001010111"; --57
            when "1001001001" => bcd_out <= "010101110001"; --571
            when "1001001010" => bcd_out <= "010101110010"; --572
            when "1001001011" => bcd_out <= "010101110011"; --573
            when "1001001100" => bcd_out <= "010101110100"; --574
            when "1001001101" => bcd_out <= "010101110101"; --575
            when "1001001110" => bcd_out <= "010101110110"; --576
            when "1001001111" => bcd_out <= "010101110111"; --577
            when "1001010000" => bcd_out <= "010101111000"; --578
            when "1001010001" => bcd_out <= "010101111001"; --579
            when "1001010010" => bcd_out <= "000001011000"; --58
            when "1001010011" => bcd_out <= "010110000001"; --581
            when "1001010100" => bcd_out <= "010110000010"; --582
            when "1001010101" => bcd_out <= "010110000011"; --583
            when "1001010110" => bcd_out <= "010110000100"; --584
            when "1001010111" => bcd_out <= "010110000101"; --585
            when "1001011000" => bcd_out <= "010110000110"; --586
            when "1001011001" => bcd_out <= "010110000111"; --587
            when "1001011010" => bcd_out <= "010110001000"; --588
            when "1001011011" => bcd_out <= "010110001001"; --589
            when "1001011100" => bcd_out <= "000001011001"; --59
            when "1001011101" => bcd_out <= "010110010001"; --591
            when "1001011110" => bcd_out <= "010110010010"; --592
            when "1001011111" => bcd_out <= "010110010011"; --593
            when "1001100000" => bcd_out <= "010110010100"; --594
            when "1001100001" => bcd_out <= "010110010101"; --595
            when "1001100010" => bcd_out <= "010110010110"; --596
            when "1001100011" => bcd_out <= "010110010111"; --597
            when "1001100100" => bcd_out <= "010110011000"; --598
            when "1001100101" => bcd_out <= "010110011001"; --599
            when "1001100110" => bcd_out <= "000000000110"; --6
            when "1001100111" => bcd_out <= "011000000001"; --601
            when "1001101000" => bcd_out <= "011000000010"; --602
            when "1001101001" => bcd_out <= "011000000011"; --603
            when "1001101010" => bcd_out <= "011000000100"; --604
            when "1001101011" => bcd_out <= "011000000100"; --604
            when "1001101100" => bcd_out <= "011000000101"; --605
            when "1001101101" => bcd_out <= "011000000110"; --606
            when "1001101110" => bcd_out <= "011000000111"; --607
            when "1001101111" => bcd_out <= "011000001000"; --608
            when "1001110000" => bcd_out <= "011000001001"; --609
            when "1001110001" => bcd_out <= "000001100001"; --61
            when "1001110010" => bcd_out <= "011000010001"; --611
            when "1001110011" => bcd_out <= "011000010010"; --612
            when "1001110100" => bcd_out <= "011000010011"; --613
            when "1001110101" => bcd_out <= "011000010100"; --614
            when "1001110110" => bcd_out <= "011000010101"; --615
            when "1001110111" => bcd_out <= "011000010110"; --616
            when "1001111000" => bcd_out <= "011000010111"; --617
            when "1001111001" => bcd_out <= "011000011000"; --618
            when "1001111010" => bcd_out <= "011000011001"; --619
            when "1001111011" => bcd_out <= "000001100010"; --62
            when "1001111100" => bcd_out <= "011000100001"; --621
            when "1001111101" => bcd_out <= "011000100010"; --622
            when "1001111110" => bcd_out <= "011000100011"; --623
            when "1001111111" => bcd_out <= "011000100100"; --624
            when "1010000000" => bcd_out <= "011000100101"; --625
            when "1010000001" => bcd_out <= "011000100110"; --626
            when "1010000010" => bcd_out <= "011000100111"; --627
            when "1010000011" => bcd_out <= "011000101000"; --628
            when "1010000100" => bcd_out <= "011000101001"; --629
            when "1010000101" => bcd_out <= "000001100011"; --63
            when "1010000110" => bcd_out <= "011000110001"; --631
            when "1010000111" => bcd_out <= "011000110010"; --632
            when "1010001000" => bcd_out <= "011000110011"; --633
            when "1010001001" => bcd_out <= "011000110100"; --634
            when "1010001010" => bcd_out <= "011000110101"; --635
            when "1010001011" => bcd_out <= "011000110110"; --636
            when "1010001100" => bcd_out <= "011000110111"; --637
            when "1010001101" => bcd_out <= "011000111000"; --638
            when "1010001110" => bcd_out <= "011000111001"; --639
            when "1010001111" => bcd_out <= "000001100100"; --64
            when "1010010000" => bcd_out <= "011001000001"; --641
            when "1010010001" => bcd_out <= "011001000010"; --642
            when "1010010010" => bcd_out <= "011001000011"; --643
            when "1010010011" => bcd_out <= "011001000100"; --644
            when "1010010100" => bcd_out <= "011001000101"; --645
            when "1010010101" => bcd_out <= "011001000110"; --646
            when "1010010110" => bcd_out <= "011001000110"; --646
            when "1010010111" => bcd_out <= "011001000111"; --647
            when "1010011000" => bcd_out <= "011001001000"; --648
            when "1010011001" => bcd_out <= "011001001001"; --649
            when "1010011010" => bcd_out <= "000001100101"; --65
            when "1010011011" => bcd_out <= "011001010001"; --651
            when "1010011100" => bcd_out <= "011001010010"; --652
            when "1010011101" => bcd_out <= "011001010011"; --653
            when "1010011110" => bcd_out <= "011001010100"; --654
            when "1010011111" => bcd_out <= "011001010101"; --655
            when "1010100000" => bcd_out <= "011001010110"; --656
            when "1010100001" => bcd_out <= "011001010111"; --657
            when "1010100010" => bcd_out <= "011001011000"; --658
            when "1010100011" => bcd_out <= "011001011001"; --659
            when "1010100100" => bcd_out <= "000001100110"; --66
            when "1010100101" => bcd_out <= "011001100001"; --661
            when "1010100110" => bcd_out <= "011001100010"; --662
            when "1010100111" => bcd_out <= "011001100011"; --663
            when "1010101000" => bcd_out <= "011001100100"; --664
            when "1010101001" => bcd_out <= "011001100101"; --665
            when "1010101010" => bcd_out <= "011001100110"; --666
            when "1010101011" => bcd_out <= "011001100111"; --667
            when "1010101100" => bcd_out <= "011001101000"; --668
            when "1010101101" => bcd_out <= "011001101001"; --669
            when "1010101110" => bcd_out <= "000001100111"; --67
            when "1010101111" => bcd_out <= "011001110001"; --671
            when "1010110000" => bcd_out <= "011001110010"; --672
            when "1010110001" => bcd_out <= "011001110011"; --673
            when "1010110010" => bcd_out <= "011001110100"; --674
            when "1010110011" => bcd_out <= "011001110101"; --675
            when "1010110100" => bcd_out <= "011001110110"; --676
            when "1010110101" => bcd_out <= "011001110111"; --677
            when "1010110110" => bcd_out <= "011001111000"; --678
            when "1010110111" => bcd_out <= "011001111001"; --679
            when "1010111000" => bcd_out <= "000001101000"; --68
            when "1010111001" => bcd_out <= "011010000001"; --681
            when "1010111010" => bcd_out <= "011010000010"; --682
            when "1010111011" => bcd_out <= "011010000011"; --683
            when "1010111100" => bcd_out <= "011010000100"; --684
            when "1010111101" => bcd_out <= "011010000101"; --685
            when "1010111110" => bcd_out <= "011010000110"; --686
            when "1010111111" => bcd_out <= "011010000111"; --687
            when "1011000000" => bcd_out <= "011010001000"; --688
            when "1011000001" => bcd_out <= "011010001000"; --688
            when "1011000010" => bcd_out <= "011010001001"; --689
            when "1011000011" => bcd_out <= "000001101001"; --69
            when "1011000100" => bcd_out <= "011010010001"; --691
            when "1011000101" => bcd_out <= "011010010010"; --692
            when "1011000110" => bcd_out <= "011010010011"; --693
            when "1011000111" => bcd_out <= "011010010100"; --694
            when "1011001000" => bcd_out <= "011010010101"; --695
            when "1011001001" => bcd_out <= "011010010110"; --696
            when "1011001010" => bcd_out <= "011010010111"; --697
            when "1011001011" => bcd_out <= "011010011000"; --698
            when "1011001100" => bcd_out <= "011010011001"; --699
            when "1011001101" => bcd_out <= "000000000111"; --7
            when "1011001110" => bcd_out <= "011100000001"; --701
            when "1011001111" => bcd_out <= "011100000010"; --702
            when "1011010000" => bcd_out <= "011100000011"; --703
            when "1011010001" => bcd_out <= "011100000100"; --704
            when "1011010010" => bcd_out <= "011100000101"; --705
            when "1011010011" => bcd_out <= "011100000110"; --706
            when "1011010100" => bcd_out <= "011100000111"; --707
            when "1011010101" => bcd_out <= "011100001000"; --708
            when "1011010110" => bcd_out <= "011100001001"; --709
            when "1011010111" => bcd_out <= "000001110001"; --71
            when "1011011000" => bcd_out <= "011100010001"; --711
            when "1011011001" => bcd_out <= "011100010010"; --712
            when "1011011010" => bcd_out <= "011100010011"; --713
            when "1011011011" => bcd_out <= "011100010100"; --714
            when "1011011100" => bcd_out <= "011100010101"; --715
            when "1011011101" => bcd_out <= "011100010110"; --716
            when "1011011110" => bcd_out <= "011100010111"; --717
            when "1011011111" => bcd_out <= "011100011000"; --718
            when "1011100000" => bcd_out <= "011100011001"; --719
            when "1011100001" => bcd_out <= "000001110010"; --72
            when "1011100010" => bcd_out <= "011100100001"; --721
            when "1011100011" => bcd_out <= "011100100010"; --722
            when "1011100100" => bcd_out <= "011100100011"; --723
            when "1011100101" => bcd_out <= "011100100100"; --724
            when "1011100110" => bcd_out <= "011100100101"; --725
            when "1011100111" => bcd_out <= "011100100110"; --726
            when "1011101000" => bcd_out <= "011100100111"; --727
            when "1011101001" => bcd_out <= "011100101000"; --728
            when "1011101010" => bcd_out <= "011100101001"; --729
            when "1011101011" => bcd_out <= "011100101001"; --729
            when "1011101100" => bcd_out <= "000001110011"; --73
            when "1011101101" => bcd_out <= "011100110001"; --731
            when "1011101110" => bcd_out <= "011100110010"; --732
            when "1011101111" => bcd_out <= "011100110011"; --733
            when "1011110000" => bcd_out <= "011100110100"; --734
            when "1011110001" => bcd_out <= "011100110101"; --735
            when "1011110010" => bcd_out <= "011100110110"; --736
            when "1011110011" => bcd_out <= "011100110111"; --737
            when "1011110100" => bcd_out <= "011100111000"; --738
            when "1011110101" => bcd_out <= "011100111001"; --739
            when "1011110110" => bcd_out <= "000001110100"; --74
            when "1011110111" => bcd_out <= "011101000001"; --741
            when "1011111000" => bcd_out <= "011101000010"; --742
            when "1011111001" => bcd_out <= "011101000011"; --743
            when "1011111010" => bcd_out <= "011101000100"; --744
            when "1011111011" => bcd_out <= "011101000101"; --745
            when "1011111100" => bcd_out <= "011101000110"; --746
            when "1011111101" => bcd_out <= "011101000111"; --747
            when "1011111110" => bcd_out <= "011101001000"; --748
            when "1011111111" => bcd_out <= "011101001001"; --749
            when "1100000000" => bcd_out <= "000001110101"; --75
            when "1100000001" => bcd_out <= "011101010001"; --751
            when "1100000010" => bcd_out <= "011101010010"; --752
            when "1100000011" => bcd_out <= "011101010011"; --753
            when "1100000100" => bcd_out <= "011101010100"; --754
            when "1100000101" => bcd_out <= "011101010101"; --755
            when "1100000110" => bcd_out <= "011101010110"; --756
            when "1100000111" => bcd_out <= "011101010111"; --757
            when "1100001000" => bcd_out <= "011101011000"; --758
            when "1100001001" => bcd_out <= "011101011001"; --759
            when "1100001010" => bcd_out <= "000001110110"; --76
            when "1100001011" => bcd_out <= "011101100001"; --761
            when "1100001100" => bcd_out <= "011101100010"; --762
            when "1100001101" => bcd_out <= "011101100011"; --763
            when "1100001110" => bcd_out <= "011101100100"; --764
            when "1100001111" => bcd_out <= "011101100101"; --765
            when "1100010000" => bcd_out <= "011101100110"; --766
            when "1100010001" => bcd_out <= "011101100111"; --767
            when "1100010010" => bcd_out <= "011101101000"; --768
            when "1100010011" => bcd_out <= "011101101001"; --769
            when "1100010100" => bcd_out <= "000001110111"; --77
            when "1100010101" => bcd_out <= "011101110001"; --771
            when "1100010110" => bcd_out <= "011101110001"; --771
            when "1100010111" => bcd_out <= "011101110010"; --772
            when "1100011000" => bcd_out <= "011101110011"; --773
            when "1100011001" => bcd_out <= "011101110100"; --774
            when "1100011010" => bcd_out <= "011101110101"; --775
            when "1100011011" => bcd_out <= "011101110110"; --776
            when "1100011100" => bcd_out <= "011101110111"; --777
            when "1100011101" => bcd_out <= "011101111000"; --778
            when "1100011110" => bcd_out <= "011101111001"; --779
            when "1100011111" => bcd_out <= "000001111000"; --78
            when "1100100000" => bcd_out <= "011110000001"; --781
            when "1100100001" => bcd_out <= "011110000010"; --782
            when "1100100010" => bcd_out <= "011110000011"; --783
            when "1100100011" => bcd_out <= "011110000100"; --784
            when "1100100100" => bcd_out <= "011110000101"; --785
            when "1100100101" => bcd_out <= "011110000110"; --786
            when "1100100110" => bcd_out <= "011110000111"; --787
            when "1100100111" => bcd_out <= "011110001000"; --788
            when "1100101000" => bcd_out <= "011110001001"; --789
            when "1100101001" => bcd_out <= "000001111001"; --79
            when "1100101010" => bcd_out <= "011110010001"; --791
            when "1100101011" => bcd_out <= "011110010010"; --792
            when "1100101100" => bcd_out <= "011110010011"; --793
            when "1100101101" => bcd_out <= "011110010100"; --794
            when "1100101110" => bcd_out <= "011110010101"; --795
            when "1100101111" => bcd_out <= "011110010110"; --796
            when "1100110000" => bcd_out <= "011110010111"; --797
            when "1100110001" => bcd_out <= "011110011000"; --798
            when "1100110010" => bcd_out <= "011110011001"; --799
            when "1100110011" => bcd_out <= "000000001000"; --8
            when "1100110100" => bcd_out <= "100000000001"; --801
            when "1100110101" => bcd_out <= "100000000010"; --802
            when "1100110110" => bcd_out <= "100000000011"; --803
            when "1100110111" => bcd_out <= "100000000100"; --804
            when "1100111000" => bcd_out <= "100000000101"; --805
            when "1100111001" => bcd_out <= "100000000110"; --806
            when "1100111010" => bcd_out <= "100000000111"; --807
            when "1100111011" => bcd_out <= "100000001000"; --808
            when "1100111100" => bcd_out <= "100000001001"; --809
            when "1100111101" => bcd_out <= "000010000001"; --81
            when "1100111110" => bcd_out <= "100000010001"; --811
            when "1100111111" => bcd_out <= "100000010010"; --812
            when "1101000000" => bcd_out <= "100000010011"; --813
            when "1101000001" => bcd_out <= "100000010011"; --813
            when "1101000010" => bcd_out <= "100000010100"; --814
            when "1101000011" => bcd_out <= "100000010101"; --815
            when "1101000100" => bcd_out <= "100000010110"; --816
            when "1101000101" => bcd_out <= "100000010111"; --817
            when "1101000110" => bcd_out <= "100000011000"; --818
            when "1101000111" => bcd_out <= "100000011001"; --819
            when "1101001000" => bcd_out <= "000010000010"; --82
            when "1101001001" => bcd_out <= "100000100001"; --821
            when "1101001010" => bcd_out <= "100000100010"; --822
            when "1101001011" => bcd_out <= "100000100011"; --823
            when "1101001100" => bcd_out <= "100000100100"; --824
            when "1101001101" => bcd_out <= "100000100101"; --825
            when "1101001110" => bcd_out <= "100000100110"; --826
            when "1101001111" => bcd_out <= "100000100111"; --827
            when "1101010000" => bcd_out <= "100000101000"; --828
            when "1101010001" => bcd_out <= "100000101001"; --829
            when "1101010010" => bcd_out <= "000010000011"; --83
            when "1101010011" => bcd_out <= "100000110001"; --831
            when "1101010100" => bcd_out <= "100000110010"; --832
            when "1101010101" => bcd_out <= "100000110011"; --833
            when "1101010110" => bcd_out <= "100000110100"; --834
            when "1101010111" => bcd_out <= "100000110101"; --835
            when "1101011000" => bcd_out <= "100000110110"; --836
            when "1101011001" => bcd_out <= "100000110111"; --837
            when "1101011010" => bcd_out <= "100000111000"; --838
            when "1101011011" => bcd_out <= "100000111001"; --839
            when "1101011100" => bcd_out <= "000010000100"; --84
            when "1101011101" => bcd_out <= "100001000001"; --841
            when "1101011110" => bcd_out <= "100001000010"; --842
            when "1101011111" => bcd_out <= "100001000011"; --843
            when "1101100000" => bcd_out <= "100001000100"; --844
            when "1101100001" => bcd_out <= "100001000101"; --845
            when "1101100010" => bcd_out <= "100001000110"; --846
            when "1101100011" => bcd_out <= "100001000111"; --847
            when "1101100100" => bcd_out <= "100001001000"; --848
            when "1101100101" => bcd_out <= "100001001001"; --849
            when "1101100110" => bcd_out <= "000010000101"; --85
            when "1101100111" => bcd_out <= "100001010001"; --851
            when "1101101000" => bcd_out <= "100001010010"; --852
            when "1101101001" => bcd_out <= "100001010011"; --853
            when "1101101010" => bcd_out <= "100001010100"; --854
            when "1101101011" => bcd_out <= "100001010100"; --854
            when "1101101100" => bcd_out <= "100001010101"; --855
            when "1101101101" => bcd_out <= "100001010110"; --856
            when "1101101110" => bcd_out <= "100001010111"; --857
            when "1101101111" => bcd_out <= "100001011000"; --858
            when "1101110000" => bcd_out <= "100001011001"; --859
            when "1101110001" => bcd_out <= "000010000110"; --86
            when "1101110010" => bcd_out <= "100001100001"; --861
            when "1101110011" => bcd_out <= "100001100010"; --862
            when "1101110100" => bcd_out <= "100001100011"; --863
            when "1101110101" => bcd_out <= "100001100100"; --864
            when "1101110110" => bcd_out <= "100001100101"; --865
            when "1101110111" => bcd_out <= "100001100110"; --866
            when "1101111000" => bcd_out <= "100001100111"; --867
            when "1101111001" => bcd_out <= "100001101000"; --868
            when "1101111010" => bcd_out <= "100001101001"; --869
            when "1101111011" => bcd_out <= "000010000111"; --87
            when "1101111100" => bcd_out <= "100001110001"; --871
            when "1101111101" => bcd_out <= "100001110010"; --872
            when "1101111110" => bcd_out <= "100001110011"; --873
            when "1101111111" => bcd_out <= "100001110100"; --874
            when "1110000000" => bcd_out <= "100001110101"; --875
            when "1110000001" => bcd_out <= "100001110110"; --876
            when "1110000010" => bcd_out <= "100001110111"; --877
            when "1110000011" => bcd_out <= "100001111000"; --878
            when "1110000100" => bcd_out <= "100001111001"; --879
            when "1110000101" => bcd_out <= "000010001000"; --88
            when "1110000110" => bcd_out <= "100010000001"; --881
            when "1110000111" => bcd_out <= "100010000010"; --882
            when "1110001000" => bcd_out <= "100010000011"; --883
            when "1110001001" => bcd_out <= "100010000100"; --884
            when "1110001010" => bcd_out <= "100010000101"; --885
            when "1110001011" => bcd_out <= "100010000110"; --886
            when "1110001100" => bcd_out <= "100010000111"; --887
            when "1110001101" => bcd_out <= "100010001000"; --888
            when "1110001110" => bcd_out <= "100010001001"; --889
            when "1110001111" => bcd_out <= "000010001001"; --89
            when "1110010000" => bcd_out <= "100010010001"; --891
            when "1110010001" => bcd_out <= "100010010010"; --892
            when "1110010010" => bcd_out <= "100010010011"; --893
            when "1110010011" => bcd_out <= "100010010100"; --894
            when "1110010100" => bcd_out <= "100010010101"; --895
            when "1110010101" => bcd_out <= "100010010110"; --896
            when "1110010110" => bcd_out <= "100010010110"; --896
            when "1110010111" => bcd_out <= "100010010111"; --897
            when "1110011000" => bcd_out <= "100010011000"; --898
            when "1110011001" => bcd_out <= "100010011001"; --899
            when "1110011010" => bcd_out <= "000000001001"; --9
            when "1110011011" => bcd_out <= "100100000001"; --901
            when "1110011100" => bcd_out <= "100100000010"; --902
            when "1110011101" => bcd_out <= "100100000011"; --903
            when "1110011110" => bcd_out <= "100100000100"; --904
            when "1110011111" => bcd_out <= "100100000101"; --905
            when "1110100000" => bcd_out <= "100100000110"; --906
            when "1110100001" => bcd_out <= "100100000111"; --907
            when "1110100010" => bcd_out <= "100100001000"; --908
            when "1110100011" => bcd_out <= "100100001001"; --909
            when "1110100100" => bcd_out <= "000010010001"; --91
            when "1110100101" => bcd_out <= "100100010001"; --911
            when "1110100110" => bcd_out <= "100100010010"; --912
            when "1110100111" => bcd_out <= "100100010011"; --913
            when "1110101000" => bcd_out <= "100100010100"; --914
            when "1110101001" => bcd_out <= "100100010101"; --915
            when "1110101010" => bcd_out <= "100100010110"; --916
            when "1110101011" => bcd_out <= "100100010111"; --917
            when "1110101100" => bcd_out <= "100100011000"; --918
            when "1110101101" => bcd_out <= "100100011001"; --919
            when "1110101110" => bcd_out <= "000010010010"; --92
            when "1110101111" => bcd_out <= "100100100001"; --921
            when "1110110000" => bcd_out <= "100100100010"; --922
            when "1110110001" => bcd_out <= "100100100011"; --923
            when "1110110010" => bcd_out <= "100100100100"; --924
            when "1110110011" => bcd_out <= "100100100101"; --925
            when "1110110100" => bcd_out <= "100100100110"; --926
            when "1110110101" => bcd_out <= "100100100111"; --927
            when "1110110110" => bcd_out <= "100100101000"; --928
            when "1110110111" => bcd_out <= "100100101001"; --929
            when "1110111000" => bcd_out <= "000010010011"; --93
            when "1110111001" => bcd_out <= "100100110001"; --931
            when "1110111010" => bcd_out <= "100100110010"; --932
            when "1110111011" => bcd_out <= "100100110011"; --933
            when "1110111100" => bcd_out <= "100100110100"; --934
            when "1110111101" => bcd_out <= "100100110101"; --935
            when "1110111110" => bcd_out <= "100100110110"; --936
            when "1110111111" => bcd_out <= "100100110111"; --937
            when "1111000000" => bcd_out <= "100100111000"; --938
            when "1111000001" => bcd_out <= "100100111000"; --938
            when "1111000010" => bcd_out <= "100100111001"; --939
            when "1111000011" => bcd_out <= "000010010100"; --94
            when "1111000100" => bcd_out <= "100101000001"; --941
            when "1111000101" => bcd_out <= "100101000010"; --942
            when "1111000110" => bcd_out <= "100101000011"; --943
            when "1111000111" => bcd_out <= "100101000100"; --944
            when "1111001000" => bcd_out <= "100101000101"; --945
            when "1111001001" => bcd_out <= "100101000110"; --946
            when "1111001010" => bcd_out <= "100101000111"; --947
            when "1111001011" => bcd_out <= "100101001000"; --948
            when "1111001100" => bcd_out <= "100101001001"; --949
            when "1111001101" => bcd_out <= "000010010101"; --95
            when "1111001110" => bcd_out <= "100101010001"; --951
            when "1111001111" => bcd_out <= "100101010010"; --952
            when "1111010000" => bcd_out <= "100101010011"; --953
            when "1111010001" => bcd_out <= "100101010100"; --954
            when "1111010010" => bcd_out <= "100101010101"; --955
            when "1111010011" => bcd_out <= "100101010110"; --956
            when "1111010100" => bcd_out <= "100101010111"; --957
            when "1111010101" => bcd_out <= "100101011000"; --958
            when "1111010110" => bcd_out <= "100101011001"; --959
            when "1111010111" => bcd_out <= "000010010110"; --96
            when "1111011000" => bcd_out <= "100101100001"; --961
            when "1111011001" => bcd_out <= "100101100010"; --962
            when "1111011010" => bcd_out <= "100101100011"; --963
            when "1111011011" => bcd_out <= "100101100100"; --964
            when "1111011100" => bcd_out <= "100101100101"; --965
            when "1111011101" => bcd_out <= "100101100110"; --966
            when "1111011110" => bcd_out <= "100101100111"; --967
            when "1111011111" => bcd_out <= "100101101000"; --968
            when "1111100000" => bcd_out <= "100101101001"; --969
            when "1111100001" => bcd_out <= "000010010111"; --97
            when "1111100010" => bcd_out <= "100101110001"; --971
            when "1111100011" => bcd_out <= "100101110010"; --972
            when "1111100100" => bcd_out <= "100101110011"; --973
            when "1111100101" => bcd_out <= "100101110100"; --974
            when "1111100110" => bcd_out <= "100101110101"; --975
            when "1111100111" => bcd_out <= "100101110110"; --976
            when "1111101000" => bcd_out <= "100101110111"; --977
            when "1111101001" => bcd_out <= "100101111000"; --978
            when "1111101010" => bcd_out <= "100101111001"; --979
            when "1111101011" => bcd_out <= "100101111001"; --979
            when "1111101100" => bcd_out <= "000010011000"; --98
            when "1111101101" => bcd_out <= "100110000001"; --981
            when "1111101110" => bcd_out <= "100110000010"; --982
            when "1111101111" => bcd_out <= "100110000011"; --983
            when "1111110000" => bcd_out <= "100110000100"; --984
            when "1111110001" => bcd_out <= "100110000101"; --985
            when "1111110010" => bcd_out <= "100110000110"; --986
            when "1111110011" => bcd_out <= "100110000111"; --987
            when "1111110100" => bcd_out <= "100110001000"; --988
            when "1111110101" => bcd_out <= "100110001001"; --989
            when "1111110110" => bcd_out <= "000010011001"; --99
            when "1111110111" => bcd_out <= "100110010001"; --991
            when "1111111000" => bcd_out <= "100110010010"; --992
            when "1111111001" => bcd_out <= "100110010011"; --993
            when "1111111010" => bcd_out <= "100110010100"; --994
            when "1111111011" => bcd_out <= "100110010101"; --995
            when "1111111100" => bcd_out <= "100110010110"; --996
            when "1111111101" => bcd_out <= "100110010111"; --997
            when "1111111110" => bcd_out <= "100110011000"; --998
            when "1111111111" => bcd_out <= "100110011001"; --999
 
			when others => null;
		end case;
	end process;
end structural;
		
	